//
// KFPC-XT Chipset
// Written by kitune-san
//
module CHIPSET (
    // Bus
    input   logic           clock,
    input   logic           reset,
);

endmodule

