//
// KFPC-XT Bus_Arbiter
// Written by kitune-san
//
module BUS_ARBITER (
    // Bus
    input   logic           clock,
    input   logic           reset,
);

endmodule

